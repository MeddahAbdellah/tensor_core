module tensor_core ();
endmodule